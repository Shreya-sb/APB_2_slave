//import uvm_pkg::*;
//`include "uvm_macros.svh"

`include "APB_2interface.sv"
`include "APB_2sequence_item.sv"
`include "APB_2sequence.sv"
`include "APB_2sequencer.sv"
`include "APB_2driver.sv"
`include "APB_2monitor_1.sv"
`include "APB_2monitor_2.sv"
`include "APB_2active_agent.sv"
`include "APB_2passive_agent.sv"
`include "APB_2scoreboard.sv"
`include "APB_2environment.sv"
`include "APB_2test.sv"
